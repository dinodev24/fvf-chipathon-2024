** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf_tb_noise.sch
**.subckt fvf_tb_noise
V1 VCC GND 1.8
I0 IBIAS GND 10u
V2 VIN GND 1.25 AC 0.2
X1 VCC GND VIN VOUT IBIAS n_fvf_cell
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.control
    noise v(VOUT) V2 dec 20 1000 1e12
    save all

    set wr_vecnames
    setplot noise1
    wrdata noise_inoise_spectrum.txt inoise_spectrum
    wrdata noise_onoise_spectrum.txt onoise_spectrum
.endc

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sym # of pins=5
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sch
.subckt n_fvf_cell VCC GND VIN VOUT IBIAS
*.ipin IBIAS
*.ipin VIN
*.opin VOUT
*.iopin GND
*.iopin VCC
X1 net1 GND VIN VOUT fvf
X2 VCC IBIAS net1 cmirror
.ends


* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/fvf.sym # of pins=4
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/fvf.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf.sch
.subckt fvf Ib GND VIN VOUT
*.ipin VIN
*.opin VOUT
*.iopin GND
*.ipin Ib
XM1 VOUT Ib GND GND sky130_fd_pr__nfet_01v8 L=0.8 W=1.29 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Ib VIN VOUT VOUT sky130_fd_pr__nfet_01v8 L=0.3 W=0.59 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/cmirror.sym # of pins=3
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/cmirror.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/cmirror.sch
.subckt cmirror VCC IIN IOUT
*.ipin IIN
*.iopin VCC
*.opin IOUT
XM1 IIN IIN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=3 W=3.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 IOUT IIN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=3 W=3.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VCC
.end
