** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf_tb_ac.sch
**.subckt fvf_tb_ac
V0 VCC GND 1.8
I0 IBIAS GND 10u
V1 VIN GND 0 AC 1
X1 VCC GND VIN VOUT IBIAS n_fvf_cell
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.control
    ac dec 20 1 1e12
    save all

    set wr_vecnames
    wrdata ac_cph_vout.txt 180*cph(v(vout))/pi
    wrdata ac_db_vout.txt db(v(vout))
    wrdata ac_vout.txt v(vout)
    exit
.endc

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sym # of pins=5
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/n_fvf_cell.sch
.subckt n_fvf_cell VCC GND VIN VOUT IBIAS
*.ipin IBIAS
*.ipin VIN
*.opin VOUT
*.iopin GND
*.iopin VCC
X1 net1 GND VIN VOUT fvf
X2 VCC IBIAS net1 cmirror
.ends


* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/fvf.sym # of pins=4
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/fvf.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf.sch
.subckt fvf Ib GND VIN VOUT
*.ipin VIN
*.opin VOUT
*.iopin GND
*.ipin Ib
XM1 Ib VIN VOUT VOUT sky130_fd_pr__nfet_01v8 L=2.5 W=1.117691 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT Ib GND GND sky130_fd_pr__nfet_01v8 L=0.6 W=1.174662 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/fvf-chipathon-2024/xschem/cmirror.sym # of pins=3
** sym_path: /foss/designs/fvf-chipathon-2024/xschem/cmirror.sym
** sch_path: /foss/designs/fvf-chipathon-2024/xschem/cmirror.sch
.subckt cmirror VCC IIN IOUT
*.ipin IIN
*.iopin VCC
*.opin IOUT
XM1 IIN IIN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 IOUT IIN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends

.GLOBAL GND
.GLOBAL VCC
.end
