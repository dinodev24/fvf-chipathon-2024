** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf_tb_noise.sch
**.subckt fvf_tb_noise
V1 VCC GND 1.8
I0 IBIAS GND 2.5u
V2 VIN GND 1.8 AC 1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.control
    noise v(Vout) V2 dec 20 1000 100e9
    save all

    set wr_vecnames
    setplot noise1
    wrdata noise_inoise_spectrum.txt inoise_spectrum
    wrdata noise_onoise_spectrum.txt onoise_spectrum
    exit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VCC
.end
