** sch_path: /foss/designs/fvf-chipathon-2024/xschem/fvf_tb_tran.sch
**.subckt fvf_tb_tran
Vin VCC GND 1.8
I0 IBIAS GND 2.5u
Vin1 VIN GND pulse(0 1.8 10ns 10ns 10ns 40ns 100ns)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.control
    tran 0.1n 1u
    save all

    set wr_vecnames
    wrdata transient_vin.txt v(vin)
    wrdata transient_vout.txt v(vout)
    exit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VCC
.end
